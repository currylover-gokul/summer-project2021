	module top_module(input [64:1]a,input [48:1]key,output[64:1]b1,b2,b3,b4,b5,b6,b7,b8,b9,b10,b11,b12,b13,b14,b15,b16);
    wire [32:1]l0,r0;
	wire [32:1] p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16;
	wire [32:1] sp1,sp2,sp3,sp4,sp5,sp6,sp7,sp8,sp9,sp10,sp11,sp12,sp13,sp14,sp15,sp16;
	wire [32:1] c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16;
    wire [48:1] e1,e2,e3,e4,e5,e6,e7,e8,e9,e10,e11,e12,e13,e14,e15,e16;
	wire [48:1] f1,f2,f3,f4,f5,f6,f7,f8,f9,f10,f11,f12,f13,f14,f15,f16;
    wire [64:1]a1;
    wire [6:1]sb1,sb2,sb3,sb4,sb5,sb6,sb7,sb8;
    wire [4:1]s1,s2,s3,s4,s5,s6,s7,s8;
    wire [6:1]sb12,sb22,sb32,sb42,sb52,sb62,sb72,sb82;
    wire [4:1]s12,s22,s32,s42,s52,s62,s72,s82;
	wire [6:1]sb13,sb23,sb33,sb43,sb53,sb63,sb73,sb83;
    wire [4:1]s13,s23,s33,s43,s53,s63,s73,s83;
    wire [6:1]sb14,sb24,sb34,sb44,sb54,sb64,sb74,sb84;
    wire [4:1]s14,s24,s34,s44,s54,s64,s74,s84;
	wire [6:1]sb15,sb25,sb35,sb45,sb55,sb65,sb75,sb85;
    wire [4:1]s15,s25,s35,s45,s55,s65,s75,s85;
    wire [6:1]sb16,sb26,sb36,sb46,sb56,sb66,sb76,sb86;
    wire [4:1]s16,s26,s36,s46,s56,s66,s76,s86;
	wire [6:1]sb17,sb27,sb37,sb47,sb57,sb67,sb77,sb87;
    wire [4:1]s17,s27,s37,s47,s57,s67,s77,s87;
    wire [6:1]sb18,sb28,sb38,sb48,sb58,sb68,sb78,sb88;
    wire [4:1]s18,s28,s38,s48,s58,s68,s78,s88;
	wire [6:1]sb19,sb29,sb39,sb49,sb59,sb69,sb79,sb89;
    wire [4:1]s19,s29,s39,s49,s59,s69,s79,s89;
	wire [6:1]sb110,sb210,sb310,sb410,sb510,sb610,sb710,sb810;
    wire [4:1]s110,s210,s310,s410,s510,s610,s710,s810;
	wire [6:1]sb111,sb211,sb311,sb411,sb511,sb611,sb711,sb811;
    wire [4:1]s111,s211,s311,s411,s511,s611,s711,s811;
	wire [6:1]sb112,sb212,sb312,sb412,sb512,sb612,sb712,sb812;
    wire [4:1]s112,s212,s312,s412,s512,s612,s712,s812;
	wire [6:1]sb113,sb213,sb313,sb413,sb513,sb613,sb713,sb813;
    wire [4:1]s113,s213,s313,s413,s513,s613,s713,s813;
	wire [6:1]sb114,sb214,sb314,sb414,sb514,sb614,sb714,sb814;
    wire [4:1]s114,s214,s314,s414,s514,s614,s714,s814;
	wire [6:1]sb115,sb215,sb315,sb415,sb515,sb615,sb715,sb815;
    wire [4:1]s115,s215,s315,s415,s515,s615,s715,s815;
	wire [6:1]sb116,sb216,sb316,sb416,sb516,sb616,sb716,sb816;
    wire [4:1]s116,s216,s316,s416,s516,s616,s716,s816;
initial_permutation I(a,l0,r0);
expansion E1(r0,e1);
assign f1 = e1 ^ key;
assign sb1=f1[48:43];
assign sb2=f1[42:37];
assign sb3=f1[36:31];
assign sb4=f1[30:25];
assign sb5=f1[24:19];
assign sb6=f1[18:13];
assign sb7=f1[12:7];
assign sb8=f1[6:1];
sbox1 S1(sb1,s1);
sbox2 S2(sb2,s2);
sbox3 S3(sb3,s3);
sbox4 S4(sb4,s4);
sbox5 S5(sb5,s5);
sbox6 S6(sb6,s6);
sbox7 S7(sb7,s7);
sbox8 S8(sb8,s8);
assign sp1={s1,s2,s3,s4,s5,s6,s7,s8};
permute P1(sp1,p1);
assign c1=p1^l0;
    assign b1={r0,c1};
    expansion E2(c1,e2);
    assign f2 = e2 ^ key;
assign sb12=f2[48:43];
assign sb22=f2[42:37];
assign sb32=f2[36:31];
assign sb42=f2[30:25];
assign sb52=f2[24:19];
assign sb62=f2[18:13];
assign sb72=f2[12:7];
assign sb82=f2[6:1];
    sbox1 S12(sb12,s12);
    sbox2 S22(sb22,s22);
    sbox3 S32(sb32,s32);
    sbox4 S42(sb42,s42);
    sbox5 S52(sb52,s52);
    sbox6 S62(sb62,s62);
    sbox7 S72(sb72,s72);
    sbox8 S82(sb82,s82);
    assign sp2={s12,s22,s32,s42,s52,s62,s72,s82};
    permute P2(sp2,p2);
    assign c2=p2^r0;
    assign b2={c1,c2};
	expansion E3(c2,e3);
    assign f3 = e3 ^ key;
assign sb13=f3[48:43];
assign sb23=f3[42:37];
assign sb33=f3[36:31];
assign sb43=f3[30:25];
assign sb53=f3[24:19];
assign sb63=f3[18:13];
assign sb73=f3[12:7];
assign sb83=f3[6:1];
    sbox1 S13(sb13,s13);
    sbox2 S23(sb23,s23);
    sbox3 S33(sb33,s33);
    sbox4 S43(sb43,s43);
    sbox5 S53(sb53,s53);
    sbox6 S63(sb63,s63);
    sbox7 S73(sb73,s73);
    sbox8 S83(sb83,s83);
    assign sp3={s13,s23,s33,s43,s53,s63,s73,s83};
    permute P3(sp3,p3);
    assign c3=p3^c1;
	assign b3={c2,c3};
expansion E4(c3,e4);
    assign f4 = e4 ^ key;
assign sb14=f4[48:43];
assign sb24=f4[42:37];
assign sb34=f4[36:31];
assign sb44=f4[30:25];
assign sb54=f4[24:19];
assign sb64=f4[18:13];
assign sb74=f4[12:7];
assign sb84=f4[6:1];  
	sbox1 S14(sb14,s14);
    sbox2 S24(sb24,s24);
    sbox3 S34(sb34,s34);
    sbox4 S44(sb44,s44);
    sbox5 S54(sb54,s54);
    sbox6 S64(sb64,s64);
    sbox7 S74(sb74,s74);
    sbox8 S84(sb84,s84);
    assign sp4={s14,s24,s34,s44,s54,s64,s74,s84};
    permute P4(sp4,p4);
    assign c4=p4^c2;
	assign b4={c3,c4};
	expansion E5(c4,e5);
    assign f5 = e5 ^ key;
assign sb15=f15[48:43];
assign sb25=f5[42:37];
assign sb35=f5[36:31];
assign sb45=f5[30:25];
assign sb55=f5[24:19];
assign sb65=f5[18:13];
assign sb75=f5[12:7];
assign sb85=f5[6:1];  
	sbox1 S15(sb15,s15);
    sbox2 S25(sb25,s25);
    sbox3 S35(sb35,s35);
    sbox4 S45(sb45,s45);
    sbox5 S55(sb55,s55);
    sbox6 S65(sb65,s65);
    sbox7 S75(sb75,s75);
    sbox8 S85(sb85,s85);
    assign sp5={s15,s25,s35,s54,sb55,s65,s75,s85};
    permute P5(sp5,p5);
    assign c5=p5^c3;
	assign b5={c4,c5};	
	expansion E6(c5,e6);
    assign f6 = e6 ^ key;
assign sb16=f6[48:43];
assign sb26=f6[42:37];
assign sb36=f6[36:31];
assign sb46=f6[30:25];
assign sb56=f6[24:19];
assign sb66=f6[18:13];
assign sb76=f6[12:7];
assign sb86=f6[6:1];  
	sbox1 S16(sb16,s16);
    sbox2 S26(sb26,s26);
    sbox3 S36(sb36,s36);
    sbox4 S46(sb46,s46);
    sbox5 S56(sb56,s56);
    sbox6 S66(sb66,s66);
    sbox7 S76(sb76,s76);
    sbox8 S86(sb86,s84);
    assign sp6={s16,s26,s36,s46,s56,s66,s76,s86};
    permute P6(sp6,p6);
    assign c6=p6^c4;
	assign b6={c5,c6};	
	expansion E7(c6,e7);
    assign f7 = e7 ^ key;
assign sb17=f7[48:43];
assign sb27=f7[42:37];
assign sb37=f7[36:31];
assign sb47=f7[30:25];
assign sb57=f7[24:19];
assign sb67=f7[18:13];
assign sb77=f7[12:7];
assign sb87=f7[6:1];  
	sbox1 S17(sb17,s17);
    sbox2 S27(sb27,s27);
    sbox3 S37(sb37,s37);
    sbox4 S47(sb47,s47);
    sbox5 S57(sb57,s57);
    sbox6 S67(sb67,s67);
    sbox7 S77(sb77,s77);
    sbox8 S87(sb87,s87);
    assign sp7={s17,s27,s37,s47,s57,s67,s77,s87};
    permute P7(sp7,p7);
    assign c7=p7^c5;
	assign b7={c6,c7};
	expansion E8(c7,e8);
    assign f8 = e8 ^ key;
assign sb18=f8[48:43];
assign sb28=f8[42:37];
assign sb38=f8[36:31];
assign sb48=f8[30:25];
assign sb58=f8[24:19];
assign sb68=f8[18:13];
assign sb78=f8[12:7];
assign sb88=f8[6:1];  
	sbox1 S18(sb18,s18);
    sbox2 S28(sb28,s28);
    sbox3 S38(sb38,s38);
    sbox4 S48(sb48,s48);
    sbox5 S58(sb58,s58);
    sbox6 S68(sb68,s68);
    sbox7 S78(sb78,s78);
    sbox8 S88(sb88,s88);
    assign sp8={s18,s28,s38,s48,s58,s68,s78,s88};
    permute P8(sp8,p8);
    assign c8=p8^c6;
	assign b8={c7,c8};
	expansion E9(c8,e9);
    assign f9 = e9 ^ key;
assign sb19=f9[48:43];
assign sb29=f9[42:37];
assign sb39=f9[36:31];
assign sb49=f9[30:25];
assign sb59=f9[24:19];
assign sb69=f9[18:13];
assign sb79=f9[12:7];
assign sb89=f9[6:1];  
	sbox1 S19(sb19,s19);
    sbox2 S29(sb29,s29);
    sbox3 S39(sb39,s39);
    sbox4 S49(sb49,s49);
    sbox5 S59(sb59,s59);
    sbox6 S69(sb69,s69);
    sbox7 S79(sb79,s79);
    sbox8 S89(sb89,s89);
    assign sp9={s19,s29,s39,s49,s59,s69,s79,s89};
    permute P9(sp9,p9);
    assign c9=p9^c7;
	assign b9={c8,c9};
	expansion E10(c9,e10);
    assign f10 = e10 ^ key;
assign sb110=f10[48:43];
assign sb210=f10[42:37];
assign sb310=f10[36:31];
assign sb410=f10[30:25];
assign sb510=f10[24:19];
assign sb610=f10[18:13];
assign sb710=f10[12:7];
assign sb810=f10[6:1];  
	sbox1 S110(sb110,s110);
    sbox2 S210(sb210,s210);
    sbox3 S310(sb310,s310);
    sbox4 S410(sb410,s410);
    sbox5 S510(sb510,s510);
    sbox6 S610(sb610,s610);
    sbox7 S710(sb710,s710);
    sbox8 S810(sb810,s810);
    assign sp10={s110,s210,s310,s410,s510,s610,s710,s810};
    permute P10(sp10,p10);
    assign c10=p10^c8;
	assign b10={c9,c10};
	expansion E11(c10,e11);
    assign f11 = e11 ^ key;
assign sb111=f11[48:43];
assign sb211=f11[42:37];
assign sb311=f11[36:31];
assign sb411=f11[30:25];
assign sb511=f11[24:19];
assign sb611=f11[18:13];
assign sb711=f11[12:7];
assign sb811=f11[6:1];  
	sbox1 S111(sb111,s111);
    sbox2 S211(sb211,s211);
    sbox3 S311(sb311,s311);
    sbox4 S411(sb411,s411);
    sbox5 S511(sb511,s511);
    sbox6 S611(sb611,s611);
    sbox7 S711(sb711,s711);
    sbox8 S811(sb811,s811);
    assign sp11={s111,s211,s311,s411,s511,s611,s711,s811};
    permute P11(sp11,p11);
    assign c11=p11^c9;
	assign b11={c10,c11};
	expansion E12(c11,e12);
    assign f12 = e12 ^ key;
assign sb112=f12[48:43];
assign sb212=f12[42:37];
assign sb312=f12[36:31];
assign sb412=f12[30:25];
assign sb512=f12[24:19];
assign sb612=f12[18:13];
assign sb712=f12[12:7];
assign sb812=f12[6:1];  
	sbox1 S112(sb112,s112);
    sbox2 S212(sb212,s212);
    sbox3 S312(sb312,s312);
    sbox4 S412(sb412,s412);
    sbox5 S512(sb512,s512);
    sbox6 S612(sb612,s612);
    sbox7 S712(sb712,s712);
    sbox8 S812(sb812,s812);
    assign sp12={s112,s212,s312,s412,s512,s612,s712,s812};
    permute P12(sp12,p12);
    assign c12=p12^c10;
	assign b12={c11,c12};
	expansion E13(c12,e13);
    assign f13 = e13 ^ key;
assign sb113=f13[48:43];
assign sb213=f13[42:37];
assign sb313=f13[36:31];
assign sb413=f13[30:25];
assign sb513=f13[24:19];
assign sb613=f13[18:13];
assign sb713=f13[12:7];
assign sb813=f13[6:1];  
	sbox1 S113(sb113,s113);
    sbox2 S213(sb213,s213);
    sbox3 S313(sb313,s313);
    sbox4 S413(sb413,s413);
    sbox5 S513(sb513,s513);
    sbox6 S613(sb613,s613);
    sbox7 S713(sb713,s713);
    sbox8 S813(sb813,s813);
    assign sp13={s113,s213,s313,s413,s513,s613,s713,s813};
    permute P13(sp13,p13);
    assign c13=p13^c11;
	assign b13={c12,c13};
	expansion E14(c13,e14);
    assign f14 = e14^ key;
assign sb114=f14[48:43];
assign sb214=f14[42:37];
assign sb314=f14[36:31];
assign sb414=f14[30:25];
assign sb514=f14[24:19];
assign sb614=f14[18:13];
assign sb714=f14[12:7];
assign sb814=f14[6:1];  
	sbox1 S114(sb114,s114);
    sbox2 S214(sb214,s214);
    sbox3 S314(sb314,s314);
    sbox4 S414(sb414,s414);
    sbox5 S514(sb514,s514);
    sbox6 S614(sb614,s614);
    sbox7 S714(sb714,s714);
    sbox8 S814(sb814,s814);
    assign sp14={s114,s214,s314,s414,s514,s614,s714,s814};
    permute P14(sp14,p14);
    assign c14=p14^c12;
	assign b14={c13,c14};
	expansion E15(c14,e15);
    assign f15 = e15^ key;
assign sb115=f15[48:43];
assign sb215=f15[42:37];
assign sb315=f15[36:31];
assign sb415=f15[30:25];
assign sb515=f15[24:19];
assign sb615=f15[18:13];
assign sb715=f15[12:7];
assign sb815=f15[6:1];  
	sbox1 S115(sb115,s115);
    sbox2 S215(sb215,s215);
    sbox3 S315(sb315,s315);
    sbox4 S415(sb415,s415);
    sbox5 S515(sb515,s515);
    sbox6 S615(sb615,s615);
    sbox7 S715(sb715,s715);
    sbox8 S815(sb815,s815);
    assign sp15={s115,s215,s315,s415,s515,s615,s715,s815};
    permute P15(sp15,p15);
    assign c15=p15^c13;
	assign b15={c14,c15};
	expansion E16(c15,e16);
    assign f16 = e16^ key;
assign sb116=f16[48:43];
assign sb216=f16[42:37];
assign sb316=f16[36:31];
assign sb416=f16[30:25];
assign sb516=f16[24:19];
assign sb616=f16[18:13];
assign sb716=f16[12:7];
assign sb816=f16[6:1];  
	sbox1 S116(sb116,s116);
    sbox2 S216(sb216,s216);
    sbox3 S316(sb316,s316);
    sbox4 S416(sb416,s416);
    sbox5 S516(sb516,s516);
    sbox6 S616(sb616,s616);
    sbox7 S716(sb716,s716);
    sbox8 S816(sb816,s816);
    assign sp16={s116,s216,s316,s416,s516,s616,s716,s816};
    permute P16(sp16,p16);
    assign c16=p16^c14;
	assign b16={c15,c16};																
endmodule
module initial_permutation(
      plaintxt,
      left_out,
    right_out);
    
    input [64:1] plaintxt;
    output [32:1] left_out;
    output [32:1] right_out;
	 
	 reg [64:1] ip;
	 assign right_out= ip[32:1] ;           
	 assign left_out= ip[64:33];          
    always@(*)begin
	            ip[1]= plaintxt[58];
					ip[2]= plaintxt[50];
					ip[3]= plaintxt[42];
					ip[4]= plaintxt[34];
					ip[5]= plaintxt[26];
					ip[6]= plaintxt[18];
					ip[7]= plaintxt[10];
					ip[8]= plaintxt[2];
					ip[9]= plaintxt[60];
					ip[10]= plaintxt[52];
					ip[11]= plaintxt[44];
					
					ip[12]= plaintxt[36];
					ip[13]= plaintxt[28];
					ip[14]= plaintxt[20];
					ip[15]= plaintxt[12];
					ip[16]= plaintxt[4];
					ip[17]= plaintxt[62];
					ip[18]= plaintxt[54];
					ip[19]= plaintxt[46];
					ip[20]= plaintxt[38];
					ip[21]= plaintxt[30];
					ip[22]= plaintxt[22];
					
					ip[23]= plaintxt[14];
					ip[24]= plaintxt[6];
					ip[25]= plaintxt[64];
					ip[26]= plaintxt[56];
					ip[27]= plaintxt[48];
					ip[28]= plaintxt[40];
					ip[29]= plaintxt[32];
					ip[30]= plaintxt[24];
					ip[31]= plaintxt[16];
					ip[32]= plaintxt[8];
					
					ip[33]= plaintxt[57];
					ip[34]= plaintxt[49];
					ip[35]= plaintxt[41];
					ip[36]= plaintxt[33];
					ip[37]= plaintxt[25];
					ip[38]= plaintxt[17];
					ip[39]= plaintxt[9];
					ip[40]= plaintxt[1];
					ip[41]= plaintxt[59];
					ip[42]= plaintxt[51];
					
					ip[43]= plaintxt[43];
					ip[44]= plaintxt[35];
					ip[45]= plaintxt[27];
					ip[46]= plaintxt[19];
					ip[47]= plaintxt[11];
					ip[48]= plaintxt[3];
					ip[49]= plaintxt[61];
					ip[50]= plaintxt[53];
					ip[51]= plaintxt[45];
					ip[52]= plaintxt[37];
					
					ip[53]= plaintxt[29];
			  		ip[54]= plaintxt[21];
					ip[55]= plaintxt[13];
					ip[56]= plaintxt[5];
					ip[57]= plaintxt[63];
					ip[58]= plaintxt[55];
					ip[59]= plaintxt[47];
					ip[60]= plaintxt[39];
					ip[61]= plaintxt[31];
					ip[62]= plaintxt[23];
					ip[63]<= plaintxt[15];
					ip[64]<= plaintxt[7];							
    end
endmodule
module expansion(input [32:1] right,output reg[48:1] ouput);
	 wire [32:1] right;
	 always @ (right)
	 begin
	 
	                      ouput[1]<= right[32];
								 ouput[2]<= right[1];
								 ouput[3]<= right[2];
								 ouput[4]<= right[3];
								 ouput[5]<= right[4];
								 ouput[6]<= right[5];
								 ouput[7]<= right[4];
								 ouput[8]<= right[5];
								 ouput[9]<= right[6];
								 ouput[10]<= right[7];
								 
								 ouput[11]<= right[8];
								 ouput[12]<= right[9];
								 ouput[13]<= right[8];
								 ouput[14]<= right[9];
								 ouput[15]<= right[10];
								 ouput[16]<= right[11];
								 ouput[17]<= right[12];
								 ouput[18]<= right[13];
								 ouput[19]<= right[12];
								 ouput[20]<= right[13];
								 
								 ouput[21]<= right[14];
								 ouput[22]<= right[15];
								 ouput[23]<= right[16];
								 ouput[24]<= right[17];
								 ouput[25]<= right[16];
								 ouput[26]<= right[17];
								 ouput[27]<= right[18];
								 ouput[28]<= right[19];
								 ouput[29]<= right[20];
								 ouput[30]<= right[21];
								 
								 ouput[31]<= right[20];
								 ouput[32]<= right[21];
								 ouput[33]<= right[22];
								 ouput[34]<= right[23];
								 ouput[35]<= right[24];
								 ouput[36]<= right[25];
								 ouput[37]<= right[24];
								 ouput[38]<= right[25];
								 ouput[39]<= right[26];
								 ouput[40]<= right[27];
								 
								 ouput[41]<= right[28];
								 ouput[42]<= right[29];
								 ouput[43]<= right[28];
								 ouput[44]<= right[29];
								 ouput[45]<= right[30];
								 ouput[46]<= right[31];
								 ouput[47]<= right[32];
								 ouput[48]<= right[1];
	 
	 end
endmodule
module sbox1(input[6:1]a,output reg [4:1]b);
    wire [6:1]a1;
assign a1={a[6],a[1],a[5:2]};
    always @(*)begin
        case(a1)
6'b000000:  b <= 4'd14;             
	 6'b000001:  b <= 4'd4;             
	 6'b000010:  b <= 4'd13;            
	 6'b000011:  b <= 4'd1;             
	 6'b000100:  b <= 4'd2;             
	 6'b000101:  b <= 4'd15;             
	 6'b000110:  b <= 4'd11;             
	 6'b000111:  b <= 4'd8;             
	 6'b001000:  b <= 4'd3;             
	 6'b001001:  b <= 4'd10;             
	 6'b001010:  b <= 4'd6;             
	 6'b001011:  b <= 4'd12;             
	 6'b001100:  b <= 4'd5;             
	 6'b001101:  b <= 4'd9;             
	 6'b001110:  b <= 4'd0;             
	 6'b001111:  b <= 4'd7;             
	 6'b010000:  b <= 4'd0;             
	 6'b010001:  b <= 4'd15;             
	 6'b010010:  b <= 4'd7;             
	 6'b010011:  b <= 4'd4;             
	 6'b010100:  b <= 4'd14;             
	 6'b010101:  b <= 4'd2;             
	 6'b010110:  b <= 4'd13;             
	 6'b010111:  b <= 4'd1;             
	 6'b011000:  b <= 4'd10;             
	 6'b011001:  b <= 4'd6;             
	 6'b011010:  b <= 4'd12;             
	 6'b011011:  b <= 4'd11;             
	 6'b011100:  b <= 4'd9;             
	 6'b011101:  b <= 4'd5;             
	 6'b011110:  b <= 4'd3;             
	 6'b011111:  b <= 4'd8;             
     6'b100000:  b <= 4'd4;             
	 6'b100001:  b <= 4'd1;             
	 6'b100010:  b <= 4'd14;             
	 6'b100011:  b <= 4'd8;             
	 6'b100100:  b <= 4'd13;             
	 6'b100101:  b <= 4'd6;             
	 6'b100110:  b <= 4'd2;             
	 6'b100111:  b <= 4'd11;             
	 6'b101000:  b <= 4'd15;             
	 6'b101001:  b <= 4'd12;             
	 6'b101010:  b <= 4'd9;             
	 6'b101011:  b <= 4'd7;             
	 6'b101100:  b <= 4'd3;             
	 6'b101101:  b <= 4'd10;             
	 6'b101110:  b <= 4'd5;             
	 6'b101111:  b <= 4'd0;             
	 6'b110000:  b <= 4'd15;             
	 6'b110001:  b <= 4'd12;             
	 6'b110010:  b <= 4'd8;             
	 6'b110011:  b <= 4'd2;             
	 6'b110100:  b <= 4'd4;             
	 6'b110101:  b <= 4'd9;            
	 6'b110110:  b <= 4'd1;             
	 6'b110111:  b <= 4'd7;            
	 6'b111000:  b <= 4'd5;        
	 6'b111001:  b <= 4'd11;        
	 6'b111010:  b <= 4'd3;       
	 6'b111011:  b <= 4'd14;       
	 6'b111100:  b <= 4'd10;       
	 6'b111101:  b <= 4'd0;       
	 6'b111110:  b <= 4'd6;      
	 6'b111111:  b <= 4'd13;      
	 default:    b <= 4'd0; 		
	 endcase 			 
	 end
endmodule
module sbox2(input[6:1]a,output reg [4:1]b);
    wire [6:1] a1; 
	 assign a1 = {a[6], a[1], a[5 : 2]}; 	  	 
	 always @(*) 	  	  
	 begin  	   	    
         case (a1)             
	 6'b000000:  b <= 4'd15;             
	 6'b000001:  b <= 4'd1;             
	 6'b000010:  b <= 4'd8;
	 6'b000011:  b <= 4'd14;             
	 6'b000100:  b <= 4'd6;             
	 6'b000101:  b <= 4'd11;             
	 6'b000110:  b <= 4'd3;             
	 6'b000111:  b <= 4'd4;             
	 6'b001000:  b <= 4'd9;             
	 6'b001001:  b <= 4'd7;             
	 6'b001010:  b <= 4'd2;             
	 6'b001011:  b <= 4'd13;             
	 6'b001100:  b <= 4'd12;             
	 6'b001101:  b <= 4'd0;             
	 6'b001110:  b <= 4'd5;             
	 6'b001111:  b <= 4'd10;             
	 6'b010000:  b <= 4'd3;             
	 6'b010001:  b <= 4'd13;             
	 6'b010010:  b <= 4'd4;             
	 6'b010011:  b <= 4'd7;             
	 6'b010100:  b <= 4'd15;             
	 6'b010101:  b <= 4'd2;             
	 6'b010110:  b <= 4'd8;             
	 6'b010111:  b <= 4'd14;             
	 6'b011000:  b <= 4'd12;             
	 6'b011001:  b <= 4'd0;             
	 6'b011010:  b <= 4'd1;             
	 6'b011011:  b <= 4'd10;             
	 6'b011100:  b <= 4'd6;             
	 6'b011101:  b <= 4'd9;             
	 6'b011110:  b <= 4'd11;             
	 6'b011111:  b <= 4'd5;             
	 6'b100000:  b <= 4'd0;             
	 6'b100001:  b <= 4'd14;             
	 6'b100010:  b <= 4'd7;             
	 6'b100011:  b <= 4'd11;             
	 6'b100100:  b <= 4'd10;             
	 6'b100101:  b <= 4'd4;             
	 6'b100110:  b <= 4'd13;             
	 6'b100111:  b <= 4'd1;             
	 6'b101000:  b <= 4'd5;             
	 6'b101001:  b <= 4'd8;             
	 6'b101010:  b <= 4'd12;             
	 6'b101011:  b <= 4'd6;             
	 6'b101100:  b <= 4'd9;             
	 6'b101101:  b <= 4'd3;             
	 6'b101110:  b <= 4'd2;             
	 6'b101111:  b <= 4'd15;             
	 6'b110000:  b <= 4'd13;             
	 6'b110001:  b <= 4'd8;             
	 6'b110010:  b <= 4'd10;             
	 6'b110011:  b <= 4'd1;             
	 6'b110100:  b <= 4'd3;             
	 6'b110101:  b <= 4'd15;            
	 6'b110110:  b <= 4'd4;             
	 6'b110111:  b <= 4'd2;            
	 6'b111000:  b <= 4'd11;        
	 6'b111001:  b <= 4'd6;        
	 6'b111010:  b <= 4'd7;       
	 6'b111011:  b <= 4'd12;       
	 6'b111100:  b <= 4'd0;       
	 6'b111101:  b <= 4'd5;       
	 6'b111110:  b <= 4'd14;      
	 6'b111111:  b <= 4'd9;      
	 default:    b <= 4'd0; 		
	 endcase 			 
	 end

endmodule
module sbox3(input [6:1] Bin, output reg [4:1] BSout);
    wire [6:1] a1;
	 assign a1 = {Bin[6], Bin[1], Bin[5 : 2]}; 	  	 
	 always @(*) 	  	  
	 begin  	   	    
         case (a1)             
	 6'b000000:  BSout <= 4'd10;             
	 6'b000001:  BSout <= 4'd0;             
	 6'b000010:  BSout <= 4'd9;            
	 6'b000011:  BSout <= 4'd14;             
	 6'b000100:  BSout <= 4'd6;             
	 6'b000101:  BSout <= 4'd3;             
	 6'b000110:  BSout <= 4'd15;             
	 6'b000111:  BSout <= 4'd5;             
	 6'b001000:  BSout <= 4'd1;             
	 6'b001001:  BSout <= 4'd13;             
	 6'b001010:  BSout <= 4'd12;             
	 6'b001011:  BSout <= 4'd7;             
	 6'b001100:  BSout <= 4'd11;             
	 6'b001101:  BSout <= 4'd4;             
	 6'b001110:  BSout <= 4'd2;             
	 6'b001111:  BSout <= 4'd8;             
	 6'b010000:  BSout <= 4'd13;             
	 6'b010001:  BSout <= 4'd7;             
	 6'b010010:  BSout <= 4'd0;             
	 6'b010011:  BSout <= 4'd9;             
	 6'b010100:  BSout <= 4'd3;             
	 6'b010101:  BSout <= 4'd4;             
	 6'b010110:  BSout <= 4'd6;             
	 6'b010111:  BSout <= 4'd10;             
	 6'b011000:  BSout <= 4'd2;             
	 6'b011001:  BSout <= 4'd8;             
	 6'b011010:  BSout <= 4'd5;             
	 6'b011011:  BSout <= 4'd14;             
	 6'b011100:  BSout <= 4'd12;             
	 6'b011101:  BSout <= 4'd11;             
	 6'b011110:  BSout <= 4'd15;             
	 6'b011111:  BSout <= 4'd1;             
	 6'b100000:  BSout <= 4'd13;             
	 6'b100001:  BSout <= 4'd6;             
	 6'b100010:  BSout <= 4'd4;             
	 6'b100011:  BSout <= 4'd9;             
	 6'b100100:  BSout <= 4'd8;             
	 6'b100101:  BSout <= 4'd15;             
	 6'b100110:  BSout <= 4'd3;             
	 6'b100111:  BSout <= 4'd0;             
	 6'b101000:  BSout <= 4'd11;             
	 6'b101001:  BSout <= 4'd1;             
	 6'b101010:  BSout <= 4'd2;             
	 6'b101011:  BSout <= 4'd12;             
	 6'b101100:  BSout <= 4'd5;             
	 6'b101101:  BSout <= 4'd10;             
	 6'b101110:  BSout <= 4'd14;             
	 6'b101111:  BSout <= 4'd7;             
	 6'b110000:  BSout <= 4'd1;             
	 6'b110001:  BSout <= 4'd10;             
	 6'b110010:  BSout <= 4'd13;             
	 6'b110011:  BSout <= 4'd0;             
	 6'b110100:  BSout <= 4'd6;             
	 6'b110101:  BSout <= 4'd9;            
	 6'b110110:  BSout <= 4'd8;             
	 6'b110111:  BSout <= 4'd7;            
	 6'b111000:  BSout <= 4'd4;        
	 6'b111001:  BSout <= 4'd15;        
	 6'b111010:  BSout <= 4'd14;       
	 6'b111011:  BSout <= 4'd3;       
	 6'b111100:  BSout <= 4'd11;       
	 6'b111101:  BSout <= 4'd5;       
	 6'b111110:  BSout <= 4'd2;      
	 6'b111111:  BSout <= 4'd12;      
	 default:    BSout <= 4'd0; 		
	 endcase 			 
	 end
endmodule
module sbox4(input [6:1] Bin,
             output reg [4:1] BSout);

     
	 wire [6:1] offset;
	  assign offset = {Bin[6], Bin[1], Bin[5 : 2]}; 	  	 
	 always @(offset) 	  	  
	 begin  	   	    
	 case (offset)             
	 6'b000000:  BSout <= 4'd7;             
	 6'b000001:  BSout <= 4'd13;             
	 6'b000010:  BSout <= 4'd14;            
	 6'b000011:  BSout <= 4'd3;             
	 6'b000100:  BSout <= 4'd0;             
	 6'b000101:  BSout <= 4'd6;             
	 6'b000110:  BSout <= 4'd9;             
	 6'b000111:  BSout <= 4'd10;             
	 6'b001000:  BSout <= 4'd1;             
	 6'b001001:  BSout <= 4'd2;             
	 6'b001010:  BSout <= 4'd8;             
	 6'b001011:  BSout <= 4'd5;             
	 6'b001100:  BSout <= 4'd11;             
	 6'b001101:  BSout <= 4'd12;             
	 6'b001110:  BSout <= 4'd4;             
	 6'b001111:  BSout <= 4'd15;             
	 6'b010000:  BSout <= 4'd13;             
	 6'b010001:  BSout <= 4'd8;             
	 6'b010010:  BSout <= 4'd11;             
	 6'b010011:  BSout <= 4'd5;             
	 6'b010100:  BSout <= 4'd6;             
	 6'b010101:  BSout <= 4'd15;             
	 6'b010110:  BSout <= 4'd0;             
	 6'b010111:  BSout <= 4'd3;             
	 6'b011000:  BSout <= 4'd4;             
	 6'b011001:  BSout <= 4'd7;             
	 6'b011010:  BSout <= 4'd2;             
	 6'b011011:  BSout <= 4'd12;             
	 6'b011100:  BSout <= 4'd1;             
	 6'b011101:  BSout <= 4'd10;             
	 6'b011110:  BSout <= 4'd14;             
	 6'b011111:  BSout <= 4'd9;             
	 6'b100000:  BSout <= 4'd10;             
	 6'b100001:  BSout <= 4'd6;             
	 6'b100010:  BSout <= 4'd9;             
	 6'b100011:  BSout <= 4'd0;             
	 6'b100100:  BSout <= 4'd12;             
	 6'b100101:  BSout <= 4'd11;             
	 6'b100110:  BSout <= 4'd7;             
	 6'b100111:  BSout <= 4'd13;             
	 6'b101000:  BSout <= 4'd15;             
	 6'b101001:  BSout <= 4'd1;             
	 6'b101010:  BSout <= 4'd3;             
	 6'b101011:  BSout <= 4'd14;             
	 6'b101100:  BSout <= 4'd5;             
	 6'b101101:  BSout <= 4'd2;             
	 6'b101110:  BSout <= 4'd8;             
	 6'b101111:  BSout <= 4'd4;             
	 6'b110000:  BSout <= 4'd3;             
	 6'b110001:  BSout <= 4'd15;             
	 6'b110010:  BSout <= 4'd0;             
	 6'b110011:  BSout <= 4'd6;             
	 6'b110100:  BSout <= 4'd10;             
	 6'b110101:  BSout <= 4'd1;            
	 6'b110110:  BSout <= 4'd13;             
	 6'b110111:  BSout <= 4'd8;            
	 6'b111000:  BSout <= 4'd9;        
	 6'b111001:  BSout <= 4'd4;        
	 6'b111010:  BSout <= 4'd5;       
	 6'b111011:  BSout <= 4'd11;       
	 6'b111100:  BSout <= 4'd12;       
	 6'b111101:  BSout <= 4'd7;       
	 6'b111110:  BSout <= 4'd2;      
	 6'b111111:  BSout <= 4'd14;      
	 default:    BSout <= 4'd0; 		
	 endcase 			 
	 end
endmodule
module sbox5(
     Bin,
    BSout
    );
    input [6:1] Bin;
    output reg [4:1] BSout;
	 wire [6:1] offset;
	  assign offset = {Bin[6], Bin[1], Bin[5 : 2]}; 	  	 
	 always @(offset) 	  	  
	 begin  	   	    
	 case (offset)             
	 6'b000000:  BSout <= 4'd2;             
	 6'b000001:  BSout <= 4'd12;             
	 6'b000010:  BSout <= 4'd4;            
	 6'b000011:  BSout <= 4'd1;             
	 6'b000100:  BSout <= 4'd7;             
	 6'b000101:  BSout <= 4'd10;             
	 6'b000110:  BSout <= 4'd11;             
	 6'b000111:  BSout <= 4'd6;             
	 6'b001000:  BSout <= 4'd8;             
	 6'b001001:  BSout <= 4'd5;             
	 6'b001010:  BSout <= 4'd3;             
	 6'b001011:  BSout <= 4'd15;             
	 6'b001100:  BSout <= 4'd13;             
	 6'b001101:  BSout <= 4'd0;             
	 6'b001110:  BSout <= 4'd14;             
	 6'b001111:  BSout <= 4'd9;             
	 6'b010000:  BSout <= 4'd14;             
	 6'b010001:  BSout <= 4'd11;             
	 6'b010010:  BSout <= 4'd2;             
	 6'b010011:  BSout <= 4'd12;             
	 6'b010100:  BSout <= 4'd4;             
	 6'b010101:  BSout <= 4'd7;             
	 6'b010110:  BSout <= 4'd13;             
	 6'b010111:  BSout <= 4'd1;             
	 6'b011000:  BSout <= 4'd5;             
	 6'b011001:  BSout <= 4'd0;             
	 6'b011010:  BSout <= 4'd15;             
	 6'b011011:  BSout <= 4'd10;             
	 6'b011100:  BSout <= 4'd3;             
	 6'b011101:  BSout <= 4'd9;             
	 6'b011110:  BSout <= 4'd8;             
	 6'b011111:  BSout <= 4'd6;             
	 6'b100000:  BSout <= 4'd4;             
	 6'b100001:  BSout <= 4'd2;             
	 6'b100010:  BSout <= 4'd1;             
	 6'b100011:  BSout <= 4'd11;             
	 6'b100100:  BSout <= 4'd10;             
	 6'b100101:  BSout <= 4'd13;             
	 6'b100110:  BSout <= 4'd7;             
	 6'b100111:  BSout <= 4'd8;             
	 6'b101000:  BSout <= 4'd15;             
	 6'b101001:  BSout <= 4'd9;             
	 6'b101010:  BSout <= 4'd12;             
	 6'b101011:  BSout <= 4'd5;             
	 6'b101100:  BSout <= 4'd6;             
	 6'b101101:  BSout <= 4'd3;             
	 6'b101110:  BSout <= 4'd0;             
	 6'b101111:  BSout <= 4'd14;             
	 6'b110000:  BSout <= 4'd11;             
	 6'b110001:  BSout <= 4'd8;             
	 6'b110010:  BSout <= 4'd12;             
	 6'b110011:  BSout <= 4'd7;             
	 6'b110100:  BSout <= 4'd1;             
	 6'b110101:  BSout <= 4'd14;            
	 6'b110110:  BSout <= 4'd2;             
	 6'b110111:  BSout <= 4'd13;            
	 6'b111000:  BSout <= 4'd6;        
	 6'b111001:  BSout <= 4'd15;        
	 6'b111010:  BSout <= 4'd0;       
	 6'b111011:  BSout <= 4'd9;       
	 6'b111100:  BSout <= 4'd10;       
	 6'b111101:  BSout <= 4'd4;       
	 6'b111110:  BSout <= 4'd5;      
	 6'b111111:  BSout <= 4'd3;      
	 default:    BSout <= 4'd0; 		
	 endcase 			 
	 end
endmodule
module sbox6(
     Bin,
     BSout
    );
	 input [6:1] Bin;
    output reg [4:1] BSout;
	 wire [6:1] offset;
	 assign offset = {Bin[6], Bin[1], Bin[5 : 2]}; 	  	 
	 always @(offset) 	  	  
	 begin  	   	    
	 case (offset)             
	 6'b000000:  BSout <= 4'd12;             
	 6'b000001:  BSout <= 4'd1;             
	 6'b000010:  BSout <= 4'd10;            
	 6'b000011:  BSout <= 4'd15;             
	 6'b000100:  BSout <= 4'd9;             
	 6'b000101:  BSout <= 4'd2;             
	 6'b000110:  BSout <= 4'd6;             
	 6'b000111:  BSout <= 4'd8;             
	 6'b001000:  BSout <= 4'd0;             
	 6'b001001:  BSout <= 4'd13;             
	 6'b001010:  BSout <= 4'd3;             
	 6'b001011:  BSout <= 4'd4;             
	 6'b001100:  BSout <= 4'd14;             
	 6'b001101:  BSout <= 4'd7;             
	 6'b001110:  BSout <= 4'd5;             
	 6'b001111:  BSout <= 4'd11;             
	 6'b010000:  BSout <= 4'd10;             
	 6'b010001:  BSout <= 4'd15;             
	 6'b010010:  BSout <= 4'd4;             
	 6'b010011:  BSout <= 4'd2;             
	 6'b010100:  BSout <= 4'd7;             
	 6'b010101:  BSout <= 4'd12;             
	 6'b010110:  BSout <= 4'd9;             
	 6'b010111:  BSout <= 4'd5;             
	 6'b011000:  BSout <= 4'd6;             
	 6'b011001:  BSout <= 4'd1;             
	 6'b011010:  BSout <= 4'd13;             
	 6'b011011:  BSout <= 4'd14;             
	 6'b011100:  BSout <= 4'd0;             
	 6'b011101:  BSout <= 4'd11;             
	 6'b011110:  BSout <= 4'd3;             
	 6'b011111:  BSout <= 4'd8;             
	 6'b100000:  BSout <= 4'd9;             
	 6'b100001:  BSout <= 4'd14;             
	 6'b100010:  BSout <= 4'd15;             
	 6'b100011:  BSout <= 4'd5;             
	 6'b100100:  BSout <= 4'd2;             
	 6'b100101:  BSout <= 4'd8;             
	 6'b100110:  BSout <= 4'd12;             
	 6'b100111:  BSout <= 4'd3;             
	 6'b101000:  BSout <= 4'd7;             
	 6'b101001:  BSout <= 4'd0;             
	 6'b101010:  BSout <= 4'd4;             
	 6'b101011:  BSout <= 4'd10;             
	 6'b101100:  BSout <= 4'd1;             
	 6'b101101:  BSout <= 4'd13;             
	 6'b101110:  BSout <= 4'd11;             
	 6'b101111:  BSout <= 4'd6;             
	 6'b110000:  BSout <= 4'd4;             
	 6'b110001:  BSout <= 4'd3;             
	 6'b110010:  BSout <= 4'd2;             
	 6'b110011:  BSout <= 4'd12;             
	 6'b110100:  BSout <= 4'd9;             
	 6'b110101:  BSout <= 4'd5;            
	 6'b110110:  BSout <= 4'd15;             
	 6'b110111:  BSout <= 4'd10;            
	 6'b111000:  BSout <= 4'd11;        
	 6'b111001:  BSout <= 4'd14;        
	 6'b111010:  BSout <= 4'd1;       
	 6'b111011:  BSout <= 4'd7;       
	 6'b111100:  BSout <= 4'd6;       
	 6'b111101:  BSout <= 4'd0;       
	 6'b111110:  BSout <= 4'd8;      
	 6'b111111:  BSout <= 4'd13;      
	 default:    BSout <= 4'd0; 		
	 endcase 			 
	 end
endmodule
module permute(
     in,
     out
    );

    input [32:1] in;
    output reg [32:1] out;
	 
	 
	 always @ (in)
	 begin 
	                    
							  out[1]<=in[16];
							  out[2]<=in[7];
							  out[3]<=in[20];
							  out[4]<=in[21];
							  out[5]<=in[29];
							  out[6]<=in[12];
							  out[7]<=in[28];
							  out[8]<=in[17];
							  out[9]<=in[1];
							  out[10]<=in[15];
							  
							  out[11]<=in[23];
							  out[12]<=in[26];
							  out[13]<=in[5];
							  out[14]<=in[18];
							  out[15]<=in[31];
							  out[16]<=in[10];
							  out[17]<=in[2];
							  out[18]<=in[8];
							  out[19]<=in[24];
							  out[20]<=in[14];
							  
							  out[21]<=in[32];
							  out[22]<=in[27];
							  out[23]<=in[3];
							  out[24]<=in[9];
							  out[25]<=in[19];
							  out[26]<=in[13];
							  out[27]<=in[30];
							  out[28]<=in[6];
							  out[29]<=in[22];
							  out[30]<=in[11];
							  
							  out[31]<=in[4];
							  out[32]<=in[25];
	 
	 
	 
	 end
endmodule
module sbox7(
     Bin,
     BSout
    );

    input [6:1] Bin;
    output reg [4:1] BSout;
	  wire [6:1] offset;
	 assign offset = {Bin[6], Bin[1], Bin[5 : 2]}; 	  	 
	 always @(offset) 	  	  
	 begin  	   	    
	 case (offset)             
	 6'b000000:  BSout <= 4'd4;             
	 6'b000001:  BSout <= 4'd11;             
	 6'b000010:  BSout <= 4'd2;            
	 6'b000011:  BSout <= 4'd14;             
	 6'b000100:  BSout <= 4'd15;             
	 6'b000101:  BSout <= 4'd0;             
	 6'b000110:  BSout <= 4'd8;             
	 6'b000111:  BSout <= 4'd13;             
	 6'b001000:  BSout <= 4'd3;             
	 6'b001001:  BSout <= 4'd12;             
	 6'b001010:  BSout <= 4'd9;             
	 6'b001011:  BSout <= 4'd7;             
	 6'b001100:  BSout <= 4'd5;             
	 6'b001101:  BSout <= 4'd10;             
	 6'b001110:  BSout <= 4'd6;             
	 6'b001111:  BSout <= 4'd1;             
	 6'b010000:  BSout <= 4'd13;             
	 6'b010001:  BSout <= 4'd0;             
	 6'b010010:  BSout <= 4'd11;             
	 6'b010011:  BSout <= 4'd7;             
	 6'b010100:  BSout <= 4'd4;             
	 6'b010101:  BSout <= 4'd9;             
	 6'b010110:  BSout <= 4'd1;             
	 6'b010111:  BSout <= 4'd10;             
	 6'b011000:  BSout <= 4'd14;             
	 6'b011001:  BSout <= 4'd3;             
	 6'b011010:  BSout <= 4'd5;             
	 6'b011011:  BSout <= 4'd12;             
	 6'b011100:  BSout <= 4'd2;             
	 6'b011101:  BSout <= 4'd15;             
	 6'b011110:  BSout <= 4'd8;             
	 6'b011111:  BSout <= 4'd6;             
	 6'b100000:  BSout <= 4'd1;             
	 6'b100001:  BSout <= 4'd4;             
	 6'b100010:  BSout <= 4'd11;             
	 6'b100011:  BSout <= 4'd13;             
	 6'b100100:  BSout <= 4'd12;             
	 6'b100101:  BSout <= 4'd3;             
	 6'b100110:  BSout <= 4'd7;             
	 6'b100111:  BSout <= 4'd14;             
	 6'b101000:  BSout <= 4'd10;             
	 6'b101001:  BSout <= 4'd15;             
	 6'b101010:  BSout <= 4'd6;             
	 6'b101011:  BSout <= 4'd8;             
	 6'b101100:  BSout <= 4'd0;             
	 6'b101101:  BSout <= 4'd5;             
	 6'b101110:  BSout <= 4'd9;             
	 6'b101111:  BSout <= 4'd2;             
	 6'b110000:  BSout <= 4'd6;             
	 6'b110001:  BSout <= 4'd11;             
	 6'b110010:  BSout <= 4'd13;             
	 6'b110011:  BSout <= 4'd8;             
	 6'b110100:  BSout <= 4'd1;             
	 6'b110101:  BSout <= 4'd4;            
	 6'b110110:  BSout <= 4'd10;             
	 6'b110111:  BSout <= 4'd7;            
	 6'b111000:  BSout <= 4'd9;        
	 6'b111001:  BSout <= 4'd5;        
	 6'b111010:  BSout <= 4'd0;       
	 6'b111011:  BSout <= 4'd15;       
	 6'b111100:  BSout <= 4'd14;       
	 6'b111101:  BSout <= 4'd2;       
	 6'b111110:  BSout <= 4'd3;      
	 6'b111111:  BSout <= 4'd12;      
	 default:    BSout <= 4'd0; 		
	 endcase 			 
	 end
	 
	 
endmodule	 
module sbox8(
     Bin,
     BSout
    );
	 
	 input [6:1] Bin;
    output reg [4:1] BSout;
	 wire [6:1] offset;
	 assign offset = {Bin[6], Bin[1], Bin[5 : 2]}; 	  	 
	 always @(offset) 	  	  
	 begin  	   	    
	 case (offset)             
	 6'b000000:  BSout <= 4'd13;             
	 6'b000001:  BSout <= 4'd2;             
	 6'b000010:  BSout <= 4'd8;            
	 6'b000011:  BSout <= 4'd4;             
	 6'b000100:  BSout <= 4'd6;             
	 6'b000101:  BSout <= 4'd15;             
	 6'b000110:  BSout <= 4'd11;             
	 6'b000111:  BSout <= 4'd1;             
	 6'b001000:  BSout <= 4'd10;             
	 6'b001001:  BSout <= 4'd9;             
	 6'b001010:  BSout <= 4'd3;             
	 6'b001011:  BSout <= 4'd14;             
	 6'b001100:  BSout <= 4'd5;             
	 6'b001101:  BSout <= 4'd0;             
	 6'b001110:  BSout <= 4'd12;             
	 6'b001111:  BSout <= 4'd7;             
	 6'b010000:  BSout <= 4'd1;             
	 6'b010001:  BSout <= 4'd15;             
	 6'b010010:  BSout <= 4'd13;             
	 6'b010011:  BSout <= 4'd8;             
	 6'b010100:  BSout <= 4'd10;             
	 6'b010101:  BSout <= 4'd3;             
	 6'b010110:  BSout <= 4'd7;             
	 6'b010111:  BSout <= 4'd4;             
	 6'b011000:  BSout <= 4'd12;             
	 6'b011001:  BSout <= 4'd5;             
	 6'b011010:  BSout <= 4'd6;             
	 6'b011011:  BSout <= 4'd11;             
	 6'b011100:  BSout <= 4'd0;             
	 6'b011101:  BSout <= 4'd14;             
	 6'b011110:  BSout <= 4'd9;             
	 6'b011111:  BSout <= 4'd2;             
	 6'b100000:  BSout <= 4'd7;             
	 6'b100001:  BSout <= 4'd11;             
	 6'b100010:  BSout <= 4'd4;             
	 6'b100011:  BSout <= 4'd1;             
	 6'b100100:  BSout <= 4'd9;             
	 6'b100101:  BSout <= 4'd12;             
	 6'b100110:  BSout <= 4'd14;             
	 6'b100111:  BSout <= 4'd2;             
	 6'b101000:  BSout <= 4'd0;             
	 6'b101001:  BSout <= 4'd6;             
	 6'b101010:  BSout <= 4'd10;             
	 6'b101011:  BSout <= 4'd13;             
	 6'b101100:  BSout <= 4'd15;             
	 6'b101101:  BSout <= 4'd3;             
	 6'b101110:  BSout <= 4'd5;             
	 6'b101111:  BSout <= 4'd8;             
	 6'b110000:  BSout <= 4'd2;             
	 6'b110001:  BSout <= 4'd1;             
	 6'b110010:  BSout <= 4'd14;             
	 6'b110011:  BSout <= 4'd7;             
	 6'b110100:  BSout <= 4'd4;             
	 6'b110101:  BSout <= 4'd10;            
	 6'b110110:  BSout <= 4'd8;             
	 6'b110111:  BSout <= 4'd13;            
	 6'b111000:  BSout <= 4'd15;        
	 6'b111001:  BSout <= 4'd12;        
	 6'b111010:  BSout <= 4'd9;       
	 6'b111011:  BSout <= 4'd0;       
	 6'b111100:  BSout <= 4'd3;       
	 6'b111101:  BSout <= 4'd5;       
	 6'b111110:  BSout <= 4'd6;      
	 6'b111111:  BSout <= 4'd11;      
	 default:    BSout <= 4'd0; 		
	 endcase 			 
	 end
	 


endmodule
module testbench;
    reg[64:1]A;
    reg [48:1]B;
    wire [64:1] g1,g2,g3,g4,g5,g6,g7,g8,g9,g10,g11,g12,g13,g14,g15,g16;
    top_module testbench(A,B,g1,g2,g3,g4,g5,g6,g7,g8,g9,g10,g11,g12,g13,g14,g15,g16);
    initial begin
        A=64'b0010101000101010001010100010101000101010001010100010101000101010;
		B=48'b101010101010101010101010101010101010101010101010;
        #1 $display ("Plaintext=%b",A);
		#1 $display ("Key=%b",B);
        #1 $display ("Cipher of round1=%b",g1);
        #1 $display ("Cipher of round2=%b",g2);
        #1 $display ("Cipher of round3=%b",g3);
        #1 $display ("Cipher of round4=%b",g4);
		#1 $display ("Cipher of round5=%b",g5);
        #1 $display ("Cipher of round6=%b",g6);
		#1 $display ("Cipher of round7=%b",g7);
        #1 $display ("Cipher of round8=%b",g8);
		#1 $display ("Cipher of round9=%b",g9);
        #1 $display ("Cipher of round10=%b",g10);
		#1 $display ("Cipher of round11=%b",g11);
        #1 $display ("Cipher of round12=%b",g12);
		#1 $display ("Cipher of round13=%b",g13);
        #1 $display ("Cipher of round14=%b",g14);
		#1 $display ("Cipher of round15=%b",g15);
        #1 $display ("Cipher of round16=%b",g16);
        $stop;
    end
endmodule
